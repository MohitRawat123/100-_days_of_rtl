`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////


module sipo(si,clk,q

    );
    input logic si,clk;
    output logic[3:0] q=0;
    always @(posedge clk)
    begin
    q[3]<=si;
    q[2]<=q[3];
    q[1]<=q[2];
    q[0]<=q[1];
    end 
endmodule
